module mixColumnsE(
       input   Input,
       output  Output
);

    //mix the columns of the input

endmodule