module createRoundKey(
       input [127:0]  RK,
       output [127:0] NextRK
);

    //create a round key from the previous round key

endmodule