module shiftRowsE(
       input   Input,
       output  Output
);

    //shift rows of the input

endmodule