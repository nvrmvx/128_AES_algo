module mixColumnsE(
    input [127:0]  Input,
    output [127:0] Output
);

//mix the columns of the input
assign Output = Input;

endmodule

//input
//d4bf5d30e0b452aeb84111f11e2798e5
//expected output
//046681e5e0cb199a48f8d37a2806264c