module shiftRowsE(
       input [127:0]  Input,
       output [127:0] Output
);

    //shift rows of the input

endmodule