module createRoundKey(
       input   RK,
       output  NextRK
);

    //create a round key from the previous round key

endmodule