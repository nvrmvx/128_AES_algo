module mixColumnsE(
       input [127:0]  Input,
       output [127:0] Output
);

    //mix the columns of the input

endmodule