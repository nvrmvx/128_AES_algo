module subBytesE(
       input [127:0]  Input,
       output [127:0] Output
);

    //substitute bytes of the input (may be hardcoded)

endmodule