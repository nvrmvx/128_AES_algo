module subBytesE(
       input   Input,
       output  Output
);

    //substitute bytes of the input (may be hardcoded)

endmodule